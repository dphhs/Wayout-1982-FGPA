`ifndef PARAMS_VH
`define PARAMS_VH

    `define MAP_WIDTH   7
    `define MAP_HEIGHT  7
    `define DATA_WIDTH  8
    `define ADDR_WIDTH  10

`endif // PARAMS_VH